module bus

