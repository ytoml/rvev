module devices

pub struct Clint {
	msip     u32
	mtimecmp u64
	mtime    u64
}
