module dram

pub const (
	// 1GiB
	dram_size = u64(0x40000000)
)