module main

import cpu

fn main() {
	c := cpu.Cpu{}
	println('${c}')
}
