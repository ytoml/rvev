module bus

pub const (
	dram_base = u64(0x80000000)
)
