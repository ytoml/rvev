module devices

import dram { Dram }

pub struct Bus {
	dram Dram
	// pub mut:
}
