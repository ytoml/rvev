module devices

pub struct Virtio {}
